// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
// CREATED		"Wed Mar 08 15:04:41 2017"

module ALU_4bit(
	Cin,
	A_next_bit,
	A_next_bit1,
	A_next_bit2,
	A_next_bit3,
	A,
	B,
	FS,
	Cout,
	F
);


input wire	Cin;
input wire	A_next_bit;
input wire	A_next_bit1;
input wire	A_next_bit2;
input wire	A_next_bit3;
input wire	[3:0] A;
input wire	[3:0] B;
input wire	[4:0] FS;
output wire	Cout;
output wire	[3:0] F;

wire	[1:0] logic1_S;
wire	[1:0] logic2_S;
wire	[1:0] logic3_S;
wire	[1:0] logic_S;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_106;
wire	SYNTHESIZED_WIRE_107;
wire	SYNTHESIZED_WIRE_108;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_109;
wire	SYNTHESIZED_WIRE_110;
wire	SYNTHESIZED_WIRE_111;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_112;
wire	SYNTHESIZED_WIRE_113;
wire	SYNTHESIZED_WIRE_114;
wire	SYNTHESIZED_WIRE_115;
wire	SYNTHESIZED_WIRE_116;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_117;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_118;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_119;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_120;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_121;
wire	SYNTHESIZED_WIRE_71;
wire	SYNTHESIZED_WIRE_72;
wire	SYNTHESIZED_WIRE_73;
wire	SYNTHESIZED_WIRE_122;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	SYNTHESIZED_WIRE_123;

assign	SYNTHESIZED_WIRE_0 = 0;
assign	SYNTHESIZED_WIRE_1 = 1;
assign	SYNTHESIZED_WIRE_3 = 0;
assign	SYNTHESIZED_WIRE_4 = 1;
assign	SYNTHESIZED_WIRE_17 = 0;
assign	SYNTHESIZED_WIRE_18 = 1;
assign	SYNTHESIZED_WIRE_30 = 0;
assign	SYNTHESIZED_WIRE_31 = 1;




FOURtoONE_MUX	b2v_inst(
	.A(FS[0]),
	.B(FS[1]),
	.C(FS[2]),
	.D(FS[3]),
	.S(logic_S),
	.Q(SYNTHESIZED_WIRE_49));


FOURtoONE_MUX	b2v_inst1(
	.A(SYNTHESIZED_WIRE_0),
	.B(SYNTHESIZED_WIRE_1),
	.C(logic_S[0]),
	.D(SYNTHESIZED_WIRE_2),
	.S(FS[2:1]),
	.Q(SYNTHESIZED_WIRE_114));



FOURtoONE_MUX	b2v_inst11(
	.A(SYNTHESIZED_WIRE_3),
	.B(SYNTHESIZED_WIRE_4),
	.C(logic1_S[0]),
	.D(SYNTHESIZED_WIRE_5),
	.S(FS[2:1]),
	.Q(SYNTHESIZED_WIRE_108));



TWOtoONE_MUX	b2v_inst13(
	.A(logic1_S[1]),
	.B(SYNTHESIZED_WIRE_6),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_107));


TWOtoONE_MUX	b2v_inst14(
	.A(SYNTHESIZED_WIRE_106),
	.B(A_next_bit1),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_15));


CarryLookaheadAdder	b2v_inst15(
	.A(SYNTHESIZED_WIRE_107),
	.B(SYNTHESIZED_WIRE_108),
	.Cin(SYNTHESIZED_WIRE_106),
	.S(SYNTHESIZED_WIRE_14));


TWOtoONE_MUX	b2v_inst16(
	.A(SYNTHESIZED_WIRE_11),
	.B(SYNTHESIZED_WIRE_12),
	.S(FS[4]),
	.Q(F[1]));


TWOtoONE_MUX	b2v_inst17(
	.A(SYNTHESIZED_WIRE_13),
	.B(logic1_S[1]),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_109));


TWOtoONE_MUX	b2v_inst18(
	.A(SYNTHESIZED_WIRE_14),
	.B(SYNTHESIZED_WIRE_15),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_12));

assign	SYNTHESIZED_WIRE_6 =  ~logic1_S[1];


TWOtoONE_MUX	b2v_inst2(
	.A(logic_S[1]),
	.B(SYNTHESIZED_WIRE_16),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_113));

assign	SYNTHESIZED_WIRE_5 =  ~logic1_S[0];




FOURtoONE_MUX	b2v_inst23(
	.A(SYNTHESIZED_WIRE_17),
	.B(SYNTHESIZED_WIRE_18),
	.C(logic2_S[0]),
	.D(SYNTHESIZED_WIRE_19),
	.S(FS[2:1]),
	.Q(SYNTHESIZED_WIRE_111));


TWOtoONE_MUX	b2v_inst24(
	.A(logic2_S[1]),
	.B(SYNTHESIZED_WIRE_20),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_110));


TWOtoONE_MUX	b2v_inst25(
	.A(SYNTHESIZED_WIRE_109),
	.B(A_next_bit2),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_29));


CarryLookaheadAdder	b2v_inst26(
	.A(SYNTHESIZED_WIRE_110),
	.B(SYNTHESIZED_WIRE_111),
	.Cin(SYNTHESIZED_WIRE_109),
	.S(SYNTHESIZED_WIRE_28));


TWOtoONE_MUX	b2v_inst27(
	.A(SYNTHESIZED_WIRE_25),
	.B(SYNTHESIZED_WIRE_26),
	.S(FS[4]),
	.Q(F[2]));


TWOtoONE_MUX	b2v_inst28(
	.A(SYNTHESIZED_WIRE_27),
	.B(logic2_S[1]),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_112));


TWOtoONE_MUX	b2v_inst29(
	.A(SYNTHESIZED_WIRE_28),
	.B(SYNTHESIZED_WIRE_29),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_26));


TWOtoONE_MUX	b2v_inst3(
	.A(Cin),
	.B(A_next_bit),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_94));

assign	SYNTHESIZED_WIRE_20 =  ~logic2_S[1];

assign	SYNTHESIZED_WIRE_19 =  ~logic2_S[0];




FOURtoONE_MUX	b2v_inst34(
	.A(SYNTHESIZED_WIRE_30),
	.B(SYNTHESIZED_WIRE_31),
	.C(logic3_S[0]),
	.D(SYNTHESIZED_WIRE_32),
	.S(FS[2:1]),
	.Q(SYNTHESIZED_WIRE_116));


TWOtoONE_MUX	b2v_inst35(
	.A(logic3_S[1]),
	.B(SYNTHESIZED_WIRE_33),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_115));


TWOtoONE_MUX	b2v_inst36(
	.A(SYNTHESIZED_WIRE_112),
	.B(A_next_bit3),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_44));


FOURtoONE_MUX	b2v_inst37(
	.A(FS[0]),
	.B(FS[1]),
	.C(FS[2]),
	.D(FS[3]),
	.S(logic1_S),
	.Q(SYNTHESIZED_WIRE_11));


FOURtoONE_MUX	b2v_inst38(
	.A(FS[0]),
	.B(FS[1]),
	.C(FS[2]),
	.D(FS[3]),
	.S(logic2_S),
	.Q(SYNTHESIZED_WIRE_25));


FOURtoONE_MUX	b2v_inst39(
	.A(FS[0]),
	.B(FS[1]),
	.C(FS[2]),
	.D(FS[3]),
	.S(logic3_S),
	.Q(SYNTHESIZED_WIRE_40));


CarryLookaheadAdder	b2v_inst4(
	.A(SYNTHESIZED_WIRE_113),
	.B(SYNTHESIZED_WIRE_114),
	.Cin(Cin),
	.S(SYNTHESIZED_WIRE_93));


CarryLookaheadAdder	b2v_inst40(
	.A(SYNTHESIZED_WIRE_115),
	.B(SYNTHESIZED_WIRE_116),
	.Cin(SYNTHESIZED_WIRE_112),
	.S(SYNTHESIZED_WIRE_43));


TWOtoONE_MUX	b2v_inst41(
	.A(SYNTHESIZED_WIRE_40),
	.B(SYNTHESIZED_WIRE_41),
	.S(FS[4]),
	.Q(F[3]));


TWOtoONE_MUX	b2v_inst42(
	.A(SYNTHESIZED_WIRE_42),
	.B(logic3_S[1]),
	.S(FS[3]),
	.Q(Cout));


TWOtoONE_MUX	b2v_inst43(
	.A(SYNTHESIZED_WIRE_43),
	.B(SYNTHESIZED_WIRE_44),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_41));

assign	SYNTHESIZED_WIRE_33 =  ~logic3_S[1];

assign	SYNTHESIZED_WIRE_32 =  ~logic3_S[0];

assign	SYNTHESIZED_WIRE_69 = SYNTHESIZED_WIRE_117 | SYNTHESIZED_WIRE_46;



assign	SYNTHESIZED_WIRE_117 = SYNTHESIZED_WIRE_114 & SYNTHESIZED_WIRE_113;


TWOtoONE_MUX	b2v_inst5(
	.A(SYNTHESIZED_WIRE_49),
	.B(SYNTHESIZED_WIRE_50),
	.S(FS[4]),
	.Q(F[0]));

assign	SYNTHESIZED_WIRE_46 = Cin & SYNTHESIZED_WIRE_118;

assign	SYNTHESIZED_WIRE_118 = SYNTHESIZED_WIRE_113 | SYNTHESIZED_WIRE_114;

assign	SYNTHESIZED_WIRE_13 = SYNTHESIZED_WIRE_54 | SYNTHESIZED_WIRE_119 | SYNTHESIZED_WIRE_56;

assign	SYNTHESIZED_WIRE_120 = SYNTHESIZED_WIRE_107 | SYNTHESIZED_WIRE_108;

assign	SYNTHESIZED_WIRE_119 = SYNTHESIZED_WIRE_108 & SYNTHESIZED_WIRE_107;

assign	SYNTHESIZED_WIRE_56 = SYNTHESIZED_WIRE_120 & SYNTHESIZED_WIRE_117;

assign	SYNTHESIZED_WIRE_54 = SYNTHESIZED_WIRE_120 & SYNTHESIZED_WIRE_118 & Cin;

assign	SYNTHESIZED_WIRE_122 = SYNTHESIZED_WIRE_110 | SYNTHESIZED_WIRE_111;

assign	SYNTHESIZED_WIRE_121 = SYNTHESIZED_WIRE_111 & SYNTHESIZED_WIRE_110;


TWOtoONE_MUX	b2v_inst6(
	.A(SYNTHESIZED_WIRE_69),
	.B(logic_S[1]),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_106));

assign	SYNTHESIZED_WIRE_27 = SYNTHESIZED_WIRE_121 | SYNTHESIZED_WIRE_71 | SYNTHESIZED_WIRE_72 | SYNTHESIZED_WIRE_73;

assign	SYNTHESIZED_WIRE_73 = SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_119;

assign	SYNTHESIZED_WIRE_71 = SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_120 & SYNTHESIZED_WIRE_117;

assign	SYNTHESIZED_WIRE_72 = SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_120 & SYNTHESIZED_WIRE_118 & Cin;

assign	SYNTHESIZED_WIRE_123 = SYNTHESIZED_WIRE_115 | SYNTHESIZED_WIRE_116;

assign	SYNTHESIZED_WIRE_86 = SYNTHESIZED_WIRE_116 & SYNTHESIZED_WIRE_115;


or5_0	b2v_inst68(
	.IN1(SYNTHESIZED_WIRE_86),
	.IN3(SYNTHESIZED_WIRE_87),
	.IN2(SYNTHESIZED_WIRE_88),
	.IN5(SYNTHESIZED_WIRE_89),
	.IN4(SYNTHESIZED_WIRE_90),
	.OUT(SYNTHESIZED_WIRE_42));

assign	SYNTHESIZED_WIRE_88 = SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_121;


TWOtoONE_MUX	b2v_inst7(
	.A(SYNTHESIZED_WIRE_93),
	.B(SYNTHESIZED_WIRE_94),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_50));

assign	SYNTHESIZED_WIRE_87 = SYNTHESIZED_WIRE_123 & SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_119;

assign	SYNTHESIZED_WIRE_90 = SYNTHESIZED_WIRE_123 & SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_120 & SYNTHESIZED_WIRE_117;


and5_1	b2v_inst72(
	.IN3(SYNTHESIZED_WIRE_120),
	.IN2(SYNTHESIZED_WIRE_122),
	.IN1(SYNTHESIZED_WIRE_123),
	.IN5(Cin),
	.IN4(SYNTHESIZED_WIRE_118),
	.OUT(SYNTHESIZED_WIRE_89));

assign	SYNTHESIZED_WIRE_16 =  ~logic_S[1];

assign	SYNTHESIZED_WIRE_2 =  ~logic_S[0];

assign	logic1_S[1] = A[1];
assign	logic1_S[0] = B[1];
assign	logic2_S[1] = A[2];
assign	logic2_S[0] = B[2];
assign	logic3_S[1] = A[3];
assign	logic3_S[0] = B[3];
assign	logic_S[0] = B[0];
assign	logic_S[1] = A[0];

endmodule

module and5_1(IN3,IN2,IN1,IN5,IN4,OUT);
/* synthesis black_box */

input IN3;
input IN2;
input IN1;
input IN5;
input IN4;
output OUT;

endmodule

module or5_0(IN1,IN3,IN2,IN5,IN4,OUT);
/* synthesis black_box */

input IN1;
input IN3;
input IN2;
input IN5;
input IN4;
output OUT;

endmodule
