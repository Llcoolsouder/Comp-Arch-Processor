library verilog;
use verilog.vl_types.all;
entity or5_0 is
    port(
        IN1             : in     vl_logic;
        IN3             : in     vl_logic;
        IN2             : in     vl_logic;
        IN5             : in     vl_logic;
        IN4             : in     vl_logic;
        \OUT\           : out    vl_logic
    );
end or5_0;
