-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Wed Feb 08 23:53:56 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY ALU_4bit IS 
	PORT
	(
		Cin :  IN  STD_LOGIC;
		A_next_bit :  IN  STD_LOGIC;
		A_next_bit1 :  IN  STD_LOGIC;
		A_next_bit2 :  IN  STD_LOGIC;
		A_next_bit3 :  IN  STD_LOGIC;
		A :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		B :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		FS :  IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		Cout :  OUT  STD_LOGIC;
		F :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ALU_4bit;

ARCHITECTURE bdf_type OF ALU_4bit IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT and5_1
	PORT(IN3 : IN STD_LOGIC;
		 IN2 : IN STD_LOGIC;
		 IN1 : IN STD_LOGIC;
		 IN5 : IN STD_LOGIC;
		 IN4 : IN STD_LOGIC;
		 OUT : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF and5_1: COMPONENT IS true;
ATTRIBUTE noopt OF and5_1: COMPONENT IS true;

COMPONENT or5_0
	PORT(IN1 : IN STD_LOGIC;
		 IN3 : IN STD_LOGIC;
		 IN2 : IN STD_LOGIC;
		 IN5 : IN STD_LOGIC;
		 IN4 : IN STD_LOGIC;
		 OUT : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF or5_0: COMPONENT IS true;
ATTRIBUTE noopt OF or5_0: COMPONENT IS true;

COMPONENT fourtoone_mux
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 S : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 Q : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT twotoone_mux
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 S : IN STD_LOGIC;
		 Q : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT carrylookaheadadder
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 Cin : IN STD_LOGIC;
		 S : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	logic1_S :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	logic2_S :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	logic3_S :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	logic_S :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_107 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_109 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_111 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_112 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_113 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_114 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_115 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_116 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_117 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_118 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_119 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_120 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_121 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_122 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_0 <= '0';
SYNTHESIZED_WIRE_1 <= '1';
SYNTHESIZED_WIRE_3 <= '0';
SYNTHESIZED_WIRE_4 <= '1';
SYNTHESIZED_WIRE_17 <= '0';
SYNTHESIZED_WIRE_18 <= '1';
SYNTHESIZED_WIRE_30 <= '0';
SYNTHESIZED_WIRE_31 <= '1';



b2v_inst : fourtoone_mux
PORT MAP(A => FS(0),
		 B => FS(1),
		 C => FS(2),
		 D => FS(3),
		 S => logic_S,
		 Q => SYNTHESIZED_WIRE_49);


b2v_inst1 : fourtoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_0,
		 B => SYNTHESIZED_WIRE_1,
		 C => logic_S(0),
		 D => SYNTHESIZED_WIRE_2,
		 S => FS(2 DOWNTO 1),
		 Q => SYNTHESIZED_WIRE_114);



b2v_inst11 : fourtoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_3,
		 B => SYNTHESIZED_WIRE_4,
		 C => logic1_S(0),
		 D => SYNTHESIZED_WIRE_5,
		 S => FS(2 DOWNTO 1),
		 Q => SYNTHESIZED_WIRE_108);



b2v_inst13 : twotoone_mux
PORT MAP(A => logic1_S(1),
		 B => SYNTHESIZED_WIRE_6,
		 S => FS(0),
		 Q => SYNTHESIZED_WIRE_107);


b2v_inst14 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_106,
		 B => A_next_bit1,
		 S => FS(0),
		 Q => SYNTHESIZED_WIRE_15);


b2v_inst15 : carrylookaheadadder
PORT MAP(A => SYNTHESIZED_WIRE_107,
		 B => SYNTHESIZED_WIRE_108,
		 Cin => SYNTHESIZED_WIRE_106,
		 S => SYNTHESIZED_WIRE_14);


b2v_inst16 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_11,
		 B => SYNTHESIZED_WIRE_12,
		 S => FS(4),
		 Q => F(1));


b2v_inst17 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_13,
		 B => logic1_S(1),
		 S => FS(3),
		 Q => SYNTHESIZED_WIRE_109);


b2v_inst18 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_14,
		 B => SYNTHESIZED_WIRE_15,
		 S => FS(3),
		 Q => SYNTHESIZED_WIRE_12);


SYNTHESIZED_WIRE_6 <= NOT(logic1_S(1));



b2v_inst2 : twotoone_mux
PORT MAP(A => logic_S(1),
		 B => SYNTHESIZED_WIRE_16,
		 S => FS(0),
		 Q => SYNTHESIZED_WIRE_113);


SYNTHESIZED_WIRE_5 <= NOT(logic1_S(0));





b2v_inst23 : fourtoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_17,
		 B => SYNTHESIZED_WIRE_18,
		 C => logic2_S(0),
		 D => SYNTHESIZED_WIRE_19,
		 S => FS(2 DOWNTO 1),
		 Q => SYNTHESIZED_WIRE_111);


b2v_inst24 : twotoone_mux
PORT MAP(A => logic2_S(1),
		 B => SYNTHESIZED_WIRE_20,
		 S => FS(0),
		 Q => SYNTHESIZED_WIRE_110);


b2v_inst25 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_109,
		 B => A_next_bit2,
		 S => FS(0),
		 Q => SYNTHESIZED_WIRE_29);


b2v_inst26 : carrylookaheadadder
PORT MAP(A => SYNTHESIZED_WIRE_110,
		 B => SYNTHESIZED_WIRE_111,
		 Cin => SYNTHESIZED_WIRE_109,
		 S => SYNTHESIZED_WIRE_28);


b2v_inst27 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_25,
		 B => SYNTHESIZED_WIRE_26,
		 S => FS(4),
		 Q => F(2));


b2v_inst28 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_27,
		 B => logic2_S(1),
		 S => FS(3),
		 Q => SYNTHESIZED_WIRE_112);


b2v_inst29 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_28,
		 B => SYNTHESIZED_WIRE_29,
		 S => FS(3),
		 Q => SYNTHESIZED_WIRE_26);


b2v_inst3 : twotoone_mux
PORT MAP(A => Cin,
		 B => A_next_bit,
		 S => FS(0),
		 Q => SYNTHESIZED_WIRE_94);


SYNTHESIZED_WIRE_20 <= NOT(logic2_S(1));



SYNTHESIZED_WIRE_19 <= NOT(logic2_S(0));





b2v_inst34 : fourtoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_30,
		 B => SYNTHESIZED_WIRE_31,
		 C => logic3_S(0),
		 D => SYNTHESIZED_WIRE_32,
		 S => FS(2 DOWNTO 1),
		 Q => SYNTHESIZED_WIRE_116);


b2v_inst35 : twotoone_mux
PORT MAP(A => logic3_S(1),
		 B => SYNTHESIZED_WIRE_33,
		 S => FS(0),
		 Q => SYNTHESIZED_WIRE_115);


b2v_inst36 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_112,
		 B => A_next_bit3,
		 S => FS(0),
		 Q => SYNTHESIZED_WIRE_44);


b2v_inst37 : fourtoone_mux
PORT MAP(A => FS(0),
		 B => FS(1),
		 C => FS(2),
		 D => FS(3),
		 S => logic1_S,
		 Q => SYNTHESIZED_WIRE_11);


b2v_inst38 : fourtoone_mux
PORT MAP(A => FS(0),
		 B => FS(1),
		 C => FS(2),
		 D => FS(3),
		 S => logic2_S,
		 Q => SYNTHESIZED_WIRE_25);


b2v_inst39 : fourtoone_mux
PORT MAP(A => FS(0),
		 B => FS(1),
		 C => FS(2),
		 D => FS(3),
		 S => logic3_S,
		 Q => SYNTHESIZED_WIRE_40);


b2v_inst4 : carrylookaheadadder
PORT MAP(A => SYNTHESIZED_WIRE_113,
		 B => SYNTHESIZED_WIRE_114,
		 Cin => Cin,
		 S => SYNTHESIZED_WIRE_93);


b2v_inst40 : carrylookaheadadder
PORT MAP(A => SYNTHESIZED_WIRE_115,
		 B => SYNTHESIZED_WIRE_116,
		 Cin => SYNTHESIZED_WIRE_112,
		 S => SYNTHESIZED_WIRE_43);


b2v_inst41 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_40,
		 B => SYNTHESIZED_WIRE_41,
		 S => FS(4),
		 Q => F(3));


b2v_inst42 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_42,
		 B => logic3_S(1),
		 S => FS(3),
		 Q => Cout);


b2v_inst43 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_43,
		 B => SYNTHESIZED_WIRE_44,
		 S => FS(3),
		 Q => SYNTHESIZED_WIRE_41);


SYNTHESIZED_WIRE_33 <= NOT(logic3_S(1));



SYNTHESIZED_WIRE_32 <= NOT(logic3_S(0));



SYNTHESIZED_WIRE_69 <= SYNTHESIZED_WIRE_117 OR SYNTHESIZED_WIRE_46;




SYNTHESIZED_WIRE_117 <= SYNTHESIZED_WIRE_114 AND SYNTHESIZED_WIRE_113;


b2v_inst5 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_49,
		 B => SYNTHESIZED_WIRE_50,
		 S => FS(4),
		 Q => F(0));


SYNTHESIZED_WIRE_46 <= Cin AND SYNTHESIZED_WIRE_118;


SYNTHESIZED_WIRE_118 <= SYNTHESIZED_WIRE_113 OR SYNTHESIZED_WIRE_114;


SYNTHESIZED_WIRE_13 <= SYNTHESIZED_WIRE_54 OR SYNTHESIZED_WIRE_119 OR SYNTHESIZED_WIRE_56;


SYNTHESIZED_WIRE_120 <= SYNTHESIZED_WIRE_107 OR SYNTHESIZED_WIRE_108;


SYNTHESIZED_WIRE_119 <= SYNTHESIZED_WIRE_108 AND SYNTHESIZED_WIRE_107;


SYNTHESIZED_WIRE_56 <= SYNTHESIZED_WIRE_120 AND SYNTHESIZED_WIRE_117;


SYNTHESIZED_WIRE_54 <= SYNTHESIZED_WIRE_120 AND SYNTHESIZED_WIRE_118 AND Cin;


SYNTHESIZED_WIRE_122 <= SYNTHESIZED_WIRE_110 OR SYNTHESIZED_WIRE_111;


SYNTHESIZED_WIRE_121 <= SYNTHESIZED_WIRE_111 AND SYNTHESIZED_WIRE_110;


b2v_inst6 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_69,
		 B => logic_S(1),
		 S => FS(3),
		 Q => SYNTHESIZED_WIRE_106);


SYNTHESIZED_WIRE_27 <= SYNTHESIZED_WIRE_121 OR SYNTHESIZED_WIRE_71 OR SYNTHESIZED_WIRE_72 OR SYNTHESIZED_WIRE_73;


SYNTHESIZED_WIRE_73 <= SYNTHESIZED_WIRE_122 AND SYNTHESIZED_WIRE_119;


SYNTHESIZED_WIRE_71 <= SYNTHESIZED_WIRE_122 AND SYNTHESIZED_WIRE_120 AND SYNTHESIZED_WIRE_117;


SYNTHESIZED_WIRE_72 <= SYNTHESIZED_WIRE_122 AND SYNTHESIZED_WIRE_120 AND SYNTHESIZED_WIRE_118 AND Cin;


SYNTHESIZED_WIRE_123 <= SYNTHESIZED_WIRE_115 OR SYNTHESIZED_WIRE_116;


SYNTHESIZED_WIRE_86 <= SYNTHESIZED_WIRE_116 AND SYNTHESIZED_WIRE_115;


b2v_inst68 : or5_0
PORT MAP(IN1 => SYNTHESIZED_WIRE_86,
		 IN3 => SYNTHESIZED_WIRE_87,
		 IN2 => SYNTHESIZED_WIRE_88,
		 IN5 => SYNTHESIZED_WIRE_89,
		 IN4 => SYNTHESIZED_WIRE_90,
		 OUT => SYNTHESIZED_WIRE_42);


SYNTHESIZED_WIRE_88 <= SYNTHESIZED_WIRE_122 AND SYNTHESIZED_WIRE_121;


b2v_inst7 : twotoone_mux
PORT MAP(A => SYNTHESIZED_WIRE_93,
		 B => SYNTHESIZED_WIRE_94,
		 S => FS(3),
		 Q => SYNTHESIZED_WIRE_50);


SYNTHESIZED_WIRE_87 <= SYNTHESIZED_WIRE_123 AND SYNTHESIZED_WIRE_122 AND SYNTHESIZED_WIRE_119;


SYNTHESIZED_WIRE_90 <= SYNTHESIZED_WIRE_123 AND SYNTHESIZED_WIRE_122 AND SYNTHESIZED_WIRE_120 AND SYNTHESIZED_WIRE_117;


b2v_inst72 : and5_1
PORT MAP(IN3 => SYNTHESIZED_WIRE_120,
		 IN2 => SYNTHESIZED_WIRE_122,
		 IN1 => SYNTHESIZED_WIRE_123,
		 IN5 => Cin,
		 IN4 => SYNTHESIZED_WIRE_118,
		 OUT => SYNTHESIZED_WIRE_89);


SYNTHESIZED_WIRE_16 <= NOT(logic_S(1));



SYNTHESIZED_WIRE_2 <= NOT(logic_S(0));



logic1_S(1) <= A(1);
logic1_S(0) <= B(1);
logic2_S(1) <= A(2);
logic2_S(0) <= B(2);
logic3_S(1) <= A(3);
logic3_S(0) <= B(3);
logic_S(0) <= B(0);
logic_S(1) <= A(0);
END bdf_type;