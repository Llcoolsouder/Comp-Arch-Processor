library verilog;
use verilog.vl_types.all;
entity and5_1 is
    port(
        IN3             : in     vl_logic;
        IN2             : in     vl_logic;
        IN1             : in     vl_logic;
        IN5             : in     vl_logic;
        IN4             : in     vl_logic;
        \OUT\           : out    vl_logic
    );
end and5_1;
