module ALU_16bit_t;
	reg Cin;
	reg [15:0]A, B;
	reg [4:0]FS;
	wire Cout;
	wire [15:0]F;
	
	