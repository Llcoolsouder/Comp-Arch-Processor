// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
// CREATED		"Mon Apr 17 20:25:09 2017"

module ALU_4bit(
	Cin,
	A_previous_bit,
	A_next_bit,
	A,
	B,
	FS,
	Cout,
	F
);


input wire	Cin;
input wire	A_previous_bit;
input wire	A_next_bit;
input wire	[3:0] A;
input wire	[3:0] B;
input wire	[4:0] FS;
output wire	Cout;
output wire	[3:0] F;

wire	[1:0] logic1_S;
wire	[1:0] logic2_S;
wire	[1:0] logic3_S;
wire	[1:0] logic_S;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_103;
wire	SYNTHESIZED_WIRE_104;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_105;
wire	SYNTHESIZED_WIRE_106;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_107;
wire	SYNTHESIZED_WIRE_108;
wire	SYNTHESIZED_WIRE_109;
wire	SYNTHESIZED_WIRE_110;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_39;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_111;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_112;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_113;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_114;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_115;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_70;
wire	SYNTHESIZED_WIRE_116;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_85;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_117;

assign	SYNTHESIZED_WIRE_0 = 0;
assign	SYNTHESIZED_WIRE_1 = 1;
assign	SYNTHESIZED_WIRE_3 = 0;
assign	SYNTHESIZED_WIRE_4 = 1;
assign	SYNTHESIZED_WIRE_16 = 0;
assign	SYNTHESIZED_WIRE_17 = 1;
assign	SYNTHESIZED_WIRE_28 = 0;
assign	SYNTHESIZED_WIRE_29 = 1;




FOURtoONE_MUX	b2v_inst(
	.A(FS[0]),
	.B(FS[1]),
	.C(FS[2]),
	.D(FS[3]),
	.S(logic_S),
	.Q(SYNTHESIZED_WIRE_46));


FOURtoONE_MUX	b2v_inst1(
	.A(SYNTHESIZED_WIRE_0),
	.B(SYNTHESIZED_WIRE_1),
	.C(logic_S[0]),
	.D(SYNTHESIZED_WIRE_2),
	.S(FS[2:1]),
	.Q(SYNTHESIZED_WIRE_108));



FOURtoONE_MUX	b2v_inst11(
	.A(SYNTHESIZED_WIRE_3),
	.B(SYNTHESIZED_WIRE_4),
	.C(logic1_S[0]),
	.D(SYNTHESIZED_WIRE_5),
	.S(FS[2:1]),
	.Q(SYNTHESIZED_WIRE_104));



TWOtoONE_MUX	b2v_inst13(
	.A(logic1_S[1]),
	.B(SYNTHESIZED_WIRE_6),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_103));


TWOtoONE_MUX	b2v_inst14(
	.A(logic_S[1]),
	.B(logic2_S[1]),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_14));


CarryLookaheadAdder	b2v_inst15(
	.A(SYNTHESIZED_WIRE_103),
	.B(SYNTHESIZED_WIRE_104),
	.Cin(SYNTHESIZED_WIRE_9),
	.S(SYNTHESIZED_WIRE_13));


TWOtoONE_MUX	b2v_inst16(
	.A(SYNTHESIZED_WIRE_10),
	.B(SYNTHESIZED_WIRE_11),
	.S(FS[4]),
	.Q(F[1]));


TWOtoONE_MUX	b2v_inst17(
	.A(SYNTHESIZED_WIRE_12),
	.B(logic1_S[1]),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_22));


TWOtoONE_MUX	b2v_inst18(
	.A(SYNTHESIZED_WIRE_13),
	.B(SYNTHESIZED_WIRE_14),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_11));

assign	SYNTHESIZED_WIRE_6 =  ~logic1_S[1];


TWOtoONE_MUX	b2v_inst2(
	.A(logic_S[1]),
	.B(SYNTHESIZED_WIRE_15),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_107));

assign	SYNTHESIZED_WIRE_5 =  ~logic1_S[0];




FOURtoONE_MUX	b2v_inst23(
	.A(SYNTHESIZED_WIRE_16),
	.B(SYNTHESIZED_WIRE_17),
	.C(logic2_S[0]),
	.D(SYNTHESIZED_WIRE_18),
	.S(FS[2:1]),
	.Q(SYNTHESIZED_WIRE_106));


TWOtoONE_MUX	b2v_inst24(
	.A(logic2_S[1]),
	.B(SYNTHESIZED_WIRE_19),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_105));


TWOtoONE_MUX	b2v_inst25(
	.A(logic1_S[1]),
	.B(logic3_S[1]),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_27));


CarryLookaheadAdder	b2v_inst26(
	.A(SYNTHESIZED_WIRE_105),
	.B(SYNTHESIZED_WIRE_106),
	.Cin(SYNTHESIZED_WIRE_22),
	.S(SYNTHESIZED_WIRE_26));


TWOtoONE_MUX	b2v_inst27(
	.A(SYNTHESIZED_WIRE_23),
	.B(SYNTHESIZED_WIRE_24),
	.S(FS[4]),
	.Q(F[2]));


TWOtoONE_MUX	b2v_inst28(
	.A(SYNTHESIZED_WIRE_25),
	.B(logic2_S[1]),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_36));


TWOtoONE_MUX	b2v_inst29(
	.A(SYNTHESIZED_WIRE_26),
	.B(SYNTHESIZED_WIRE_27),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_24));


TWOtoONE_MUX	b2v_inst3(
	.A(A_previous_bit),
	.B(logic1_S[1]),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_91));

assign	SYNTHESIZED_WIRE_19 =  ~logic2_S[1];

assign	SYNTHESIZED_WIRE_18 =  ~logic2_S[0];




FOURtoONE_MUX	b2v_inst34(
	.A(SYNTHESIZED_WIRE_28),
	.B(SYNTHESIZED_WIRE_29),
	.C(logic3_S[0]),
	.D(SYNTHESIZED_WIRE_30),
	.S(FS[2:1]),
	.Q(SYNTHESIZED_WIRE_110));


TWOtoONE_MUX	b2v_inst35(
	.A(logic3_S[1]),
	.B(SYNTHESIZED_WIRE_31),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_109));


TWOtoONE_MUX	b2v_inst36(
	.A(logic2_S[1]),
	.B(A_next_bit),
	.S(FS[0]),
	.Q(SYNTHESIZED_WIRE_41));


FOURtoONE_MUX	b2v_inst37(
	.A(FS[0]),
	.B(FS[1]),
	.C(FS[2]),
	.D(FS[3]),
	.S(logic1_S),
	.Q(SYNTHESIZED_WIRE_10));


FOURtoONE_MUX	b2v_inst38(
	.A(FS[0]),
	.B(FS[1]),
	.C(FS[2]),
	.D(FS[3]),
	.S(logic2_S),
	.Q(SYNTHESIZED_WIRE_23));


FOURtoONE_MUX	b2v_inst39(
	.A(FS[0]),
	.B(FS[1]),
	.C(FS[2]),
	.D(FS[3]),
	.S(logic3_S),
	.Q(SYNTHESIZED_WIRE_37));


CarryLookaheadAdder	b2v_inst4(
	.A(SYNTHESIZED_WIRE_107),
	.B(SYNTHESIZED_WIRE_108),
	.Cin(Cin),
	.S(SYNTHESIZED_WIRE_90));


CarryLookaheadAdder	b2v_inst40(
	.A(SYNTHESIZED_WIRE_109),
	.B(SYNTHESIZED_WIRE_110),
	.Cin(SYNTHESIZED_WIRE_36),
	.S(SYNTHESIZED_WIRE_40));


TWOtoONE_MUX	b2v_inst41(
	.A(SYNTHESIZED_WIRE_37),
	.B(SYNTHESIZED_WIRE_38),
	.S(FS[4]),
	.Q(F[3]));


TWOtoONE_MUX	b2v_inst42(
	.A(SYNTHESIZED_WIRE_39),
	.B(logic3_S[1]),
	.S(FS[3]),
	.Q(Cout));


TWOtoONE_MUX	b2v_inst43(
	.A(SYNTHESIZED_WIRE_40),
	.B(SYNTHESIZED_WIRE_41),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_38));

assign	SYNTHESIZED_WIRE_31 =  ~logic3_S[1];

assign	SYNTHESIZED_WIRE_30 =  ~logic3_S[0];

assign	SYNTHESIZED_WIRE_66 = SYNTHESIZED_WIRE_111 | SYNTHESIZED_WIRE_43;



assign	SYNTHESIZED_WIRE_111 = SYNTHESIZED_WIRE_108 & SYNTHESIZED_WIRE_107;


TWOtoONE_MUX	b2v_inst5(
	.A(SYNTHESIZED_WIRE_46),
	.B(SYNTHESIZED_WIRE_47),
	.S(FS[4]),
	.Q(F[0]));

assign	SYNTHESIZED_WIRE_43 = Cin & SYNTHESIZED_WIRE_112;

assign	SYNTHESIZED_WIRE_112 = SYNTHESIZED_WIRE_107 | SYNTHESIZED_WIRE_108;

assign	SYNTHESIZED_WIRE_12 = SYNTHESIZED_WIRE_51 | SYNTHESIZED_WIRE_113 | SYNTHESIZED_WIRE_53;

assign	SYNTHESIZED_WIRE_114 = SYNTHESIZED_WIRE_103 | SYNTHESIZED_WIRE_104;

assign	SYNTHESIZED_WIRE_113 = SYNTHESIZED_WIRE_104 & SYNTHESIZED_WIRE_103;

assign	SYNTHESIZED_WIRE_53 = SYNTHESIZED_WIRE_114 & SYNTHESIZED_WIRE_111;

assign	SYNTHESIZED_WIRE_51 = SYNTHESIZED_WIRE_114 & SYNTHESIZED_WIRE_112 & Cin;

assign	SYNTHESIZED_WIRE_116 = SYNTHESIZED_WIRE_105 | SYNTHESIZED_WIRE_106;

assign	SYNTHESIZED_WIRE_115 = SYNTHESIZED_WIRE_106 & SYNTHESIZED_WIRE_105;


TWOtoONE_MUX	b2v_inst6(
	.A(SYNTHESIZED_WIRE_66),
	.B(logic_S[1]),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_9));

assign	SYNTHESIZED_WIRE_25 = SYNTHESIZED_WIRE_115 | SYNTHESIZED_WIRE_68 | SYNTHESIZED_WIRE_69 | SYNTHESIZED_WIRE_70;

assign	SYNTHESIZED_WIRE_70 = SYNTHESIZED_WIRE_116 & SYNTHESIZED_WIRE_113;

assign	SYNTHESIZED_WIRE_68 = SYNTHESIZED_WIRE_116 & SYNTHESIZED_WIRE_114 & SYNTHESIZED_WIRE_111;

assign	SYNTHESIZED_WIRE_69 = SYNTHESIZED_WIRE_116 & SYNTHESIZED_WIRE_114 & SYNTHESIZED_WIRE_112 & Cin;

assign	SYNTHESIZED_WIRE_117 = SYNTHESIZED_WIRE_109 | SYNTHESIZED_WIRE_110;

assign	SYNTHESIZED_WIRE_83 = SYNTHESIZED_WIRE_110 & SYNTHESIZED_WIRE_109;


or5_0	b2v_inst68(
	.IN1(SYNTHESIZED_WIRE_83),
	.IN3(SYNTHESIZED_WIRE_84),
	.IN2(SYNTHESIZED_WIRE_85),
	.IN5(SYNTHESIZED_WIRE_86),
	.IN4(SYNTHESIZED_WIRE_87),
	.OUT(SYNTHESIZED_WIRE_39));

assign	SYNTHESIZED_WIRE_85 = SYNTHESIZED_WIRE_116 & SYNTHESIZED_WIRE_115;


TWOtoONE_MUX	b2v_inst7(
	.A(SYNTHESIZED_WIRE_90),
	.B(SYNTHESIZED_WIRE_91),
	.S(FS[3]),
	.Q(SYNTHESIZED_WIRE_47));

assign	SYNTHESIZED_WIRE_84 = SYNTHESIZED_WIRE_117 & SYNTHESIZED_WIRE_116 & SYNTHESIZED_WIRE_113;

assign	SYNTHESIZED_WIRE_87 = SYNTHESIZED_WIRE_117 & SYNTHESIZED_WIRE_116 & SYNTHESIZED_WIRE_114 & SYNTHESIZED_WIRE_111;


and5_1	b2v_inst72(
	.IN3(SYNTHESIZED_WIRE_114),
	.IN2(SYNTHESIZED_WIRE_116),
	.IN1(SYNTHESIZED_WIRE_117),
	.IN5(Cin),
	.IN4(SYNTHESIZED_WIRE_112),
	.OUT(SYNTHESIZED_WIRE_86));

assign	SYNTHESIZED_WIRE_15 =  ~logic_S[1];

assign	SYNTHESIZED_WIRE_2 =  ~logic_S[0];

assign	logic1_S[0] = B[1];
assign	logic1_S[1] = A[1];
assign	logic2_S[0] = B[2];
assign	logic2_S[1] = A[2];
assign	logic3_S[0] = B[3];
assign	logic3_S[1] = A[3];
assign	logic_S[0] = B[0];
assign	logic_S[1] = A[0];

endmodule

module and5_1(IN3,IN2,IN1,IN5,IN4,OUT);
/* synthesis black_box */

input IN3;
input IN2;
input IN1;
input IN5;
input IN4;
output OUT;

endmodule

module or5_0(IN1,IN3,IN2,IN5,IN4,OUT);
/* synthesis black_box */

input IN1;
input IN3;
input IN2;
input IN5;
input IN4;
output OUT;

endmodule
