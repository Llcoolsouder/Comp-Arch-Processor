library verilog;
use verilog.vl_types.all;
entity ALU_16bit_tb is
end ALU_16bit_tb;
