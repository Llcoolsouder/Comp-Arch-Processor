library verilog;
use verilog.vl_types.all;
entity ALU_16bit_t is
end ALU_16bit_t;
