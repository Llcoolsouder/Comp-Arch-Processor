library verilog;
use verilog.vl_types.all;
entity Top_Level_ModelSim_v_t is
end Top_Level_ModelSim_v_t;
