module rom_case(out, PC);
    output reg[15:0] out;
    input [7:0] PC; //address- 8 deep memory
    
    always @(PC) begin
        case(PC)
   
        //CLR
        8'b00000000 : out[15:0]<=16'b0100000001001010;//DA=1,AA=X,BA=X
    
        //ADDI
        8'b00000001 : out[15:0]<=16'b0000100100000001;//reg 1 lit 1
        
        //SUBI
        8'b00000010 : out[15:0]<=16'b0001001000000001;//reg2 lit 1
        
        //ANDI
        8'b00000011 : out[15:0]<=16'b0001101100000001;//reg 3 lit 1
        
        //ORI
        8'b00000100 : out[15:0]<=16'b0010110000000001;//reg 4 lit 1
        
        //XORI
        8'b00000101 : out[15:0]<=16'b0011010100000001;//reg 5 lit 1
        
        //01 Operations 7 op code DA,AA,BA
        
         //INC
        8'b00000110 : out[15:0]<=16'b0110000001001000;//DA=1,AA=1,BA=X
        
        //ADD
        8'b00000111 : out[15:0]<=16'b0110100001001010;//DA=1,AA=1,BA=2
        
        //ADDC
        8'b00001000 : out[15:0]<=16'b0110101001001010;//DA=1,AA=1,BA=2
        
        //SUB
        8'b00001001 : out[15:0]<=16'b0110110001001010;//DA=1,AA=1,BA=2
        
        //DEC
        8'b00001010 : out[15:0]<=16'b0110010001001000;//DA=1,AA=1,BA=X
        
        //NEG
        8'b00001011 : out[15:0]<=16'b0110001011001000;//DA=3,AA=1,BA=X
        
        //SHR
        8'b00001100 : out[15:0]<=16'b0111001001001010;//DA=1,AA=1,BA=X
        
        //SHL
        8'b00001101 : out[15:0]<=16'b0111000001001010;//DA=1,AA=1,B=X
        
        //CLR
        8'b00001110 : out[15:0]<=16'b0100000001001010;//DA=1,AA=X,BA=X
        
        //SET
        8'b00001111 : out[15:0]<=16'b0101111001001010;//DA=1,AA=X,BA=X
        
        //NOT
        8'b00010000 :out[15:0]<=16'b0100011101001010;//DA=5,AA=1,BA=X
        
        //AND
        8'b00010001 : out[15:0]<=16'b0101000001001010;//DA=1,AA=1,BA=2
        
        //OR
        8'b00010010 : out[15:0]<=16'b0101110001001010;//DA=1,AA=1,BA=2
        
        //XOR
        8'b00010011 : out[15:0]<=16'b0100110001001010;//DA=1,AA=1,BA=2
        
        //MOVA
        8'b00010100 : out[15:0]<=16'b0101100111001010;//DA=7,AA=1,BA=X
        
        //MOVB
        8'b00010101 : out[15:0]<=16'b0101010110001010;//DA=6,AA=X,BA=2
        
        
        //10 Operations
        //LRLI(EX0)
        8'b00010110 : out[15:0]<=16'b1000010001001010;//DA=1,AA=X,BA=X
        
        //LRLI(EX1)
        8'b00010111 : out[15:0]<=16'b0000000000000001;//constant = 1
        
        //LDI
        8'b00011000 : out[15:0]<=16'b1010000100000001;//reg 1 lit 1
        
        //STI
        8'b00011001 : out[15:0]<=16'b1010101000000001;//reg2 lit 1
        
        //Push
        8'b00011010 : out[15:0]<=16'b1000000001001010;//DA=1,AA=1,BA=2
        
        //Pop
        8'b00011011 : out[15:0]<=16'b1000001001001010;//DA=1,AA=1,BA=2
        
        //STR
        8'b00011100 : out[15:0]<=16'b1000101001001010;//DA=1,AA=1,BA=2
        
        //LDR
        8'b00011101 : out[15:0]<=16'b1000100001001010;//DA=1,AA=1,BA=2
        
        //CALL(EX0)
        8'b00011110 : out[15:0]<=16'b1001110000000100;//lit = 4
        
        //RET
        8'b00011111 : out[15:0]<=16'b1001111001001010;//do not cares
        
        //BRZ
        8'b00100000 : out[15:0]<=16'b1011001100000001;//reg 3 lit 1
        
        //BRN
        8'b00100001 : out[15:0]<=16'b1011110000000001;//reg 4 lit 1
        
        //BSET
        8'b00100010 : out[15:0]<=16'b1001001001001010;//DA=1,AA=1,BA=2
        
        //BCLR
        8'b00100011 : out[15:0]<=16'b1001000001001010;//DA=1,AA=1,BA=2
        
        //JMPR
        8'b00100100 : out[15:0]<=16'b1001101001001010;//DA=1,AA=1,BA=2
        
        
        //11 Operation 2 bit op, 3bit DA, 11 bit lit
        
        8'b00100101 : out[15:0] <= 16'b1101100000000001; //DA is reg 3 and literal is d1
        default: out = 16'b0000000000000000; //NOP

        endcase
    end
endmodule // rom_case