module ALU_16bit_tb;


endmodule
	
	