library verilog;
use verilog.vl_types.all;
entity Register_File_t is
end Register_File_t;
