module address_selector(
	input [15:0]ADD,
	output  reg [16:0]Q,
	output reg RAM_S
	);
	
	always @* begin
		if (ADD[15:0]<17) begin
			RAM_S<=1'b0;
		end 
		else begin
			RAM_S<=1'b1;
		end
		case (ADD)
			16'h0000: 	Q<=17'b00000000000000001;
			16'h0001: 	Q<=17'b00000000000000010;
			16'h0002: 	Q<=17'b00000000000000100;
			16'h0003: 	Q<=17'b00000000000001000;
			16'h0004: 	Q<=17'b00000000000010000;
			16'h0005: 	Q<=17'b00000000000100000;
			16'h0006: 	Q<=17'b00000000001000000;
			16'h0007: 	Q<=17'b00000000010000000;
			16'h0008: 	Q<=17'b00000000100000000;
			16'h0009: 	Q<=17'b00000001000000000;
			16'h000a: 	Q<=17'b00000010000000000;
			16'h000b: 	Q<=17'b00000100000000000;
			16'h000c: 	Q<=17'b00001000000000000;
			16'h000d: 	Q<=17'b00010000000000000;
			16'h000e: 	Q<=17'b00100000000000000;
			16'h000f: 	Q<=17'b01000000000000000;
			16'h0010: 	Q<=17'b10000000000000000;
			default:		Q<=17'b00000000000000000;	
		endcase
	end
endmodule
			