`define LRLI
`define RET
 
module ControlUnitFSM(Instr, CLK, CW);
	input [15:0]Instr;
	input CLK;
	output reg [52:0]CW;
	
	//case (Instr)
	//	default:
	//endcase
	
endmodule 

//module ControlUnitDecoder_0 (
	
//);